VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cla
  CLASS BLOCK ;
  FOREIGN cla ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 17.360 0.000 17.920 4.000 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 0.000 50.960 4.000 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 83.440 0.000 84.000 4.000 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END A[3]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.520 0.000 150.080 4.000 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 182.560 0.000 183.120 4.000 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.600 0.000 216.160 4.000 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 0.000 249.200 4.000 ;
    END
  END B[3]
  PIN S[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 29.680 296.000 30.240 300.000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 89.600 296.000 90.160 300.000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 149.520 296.000 150.080 300.000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 209.440 296.000 210.000 300.000 ;
    END
  END S[3]
  PIN cin
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.680 0.000 282.240 4.000 ;
    END
  END cin
  PIN cout
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 269.360 296.000 269.920 300.000 ;
    END
  END cout
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 292.880 283.210 ;
      LAYER Metal2 ;
        RECT 16.380 295.700 29.380 296.000 ;
        RECT 30.540 295.700 89.300 296.000 ;
        RECT 90.460 295.700 149.220 296.000 ;
        RECT 150.380 295.700 209.140 296.000 ;
        RECT 210.300 295.700 269.060 296.000 ;
        RECT 270.220 295.700 287.140 296.000 ;
        RECT 16.380 4.300 287.140 295.700 ;
        RECT 16.380 4.000 17.060 4.300 ;
        RECT 18.220 4.000 50.100 4.300 ;
        RECT 51.260 4.000 83.140 4.300 ;
        RECT 84.300 4.000 116.180 4.300 ;
        RECT 117.340 4.000 149.220 4.300 ;
        RECT 150.380 4.000 182.260 4.300 ;
        RECT 183.420 4.000 215.300 4.300 ;
        RECT 216.460 4.000 248.340 4.300 ;
        RECT 249.500 4.000 281.380 4.300 ;
        RECT 282.540 4.000 287.140 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 15.540 287.190 282.380 ;
  END
END cla
END LIBRARY

