magic
tech gf180mcuC
magscale 1 5
timestamp 1670225163
<< obsm1 >>
rect 672 1538 29288 28321
<< metal2 >>
rect 2968 29600 3024 30000
rect 8960 29600 9016 30000
rect 14952 29600 15008 30000
rect 20944 29600 21000 30000
rect 26936 29600 26992 30000
rect 1736 0 1792 400
rect 5040 0 5096 400
rect 8344 0 8400 400
rect 11648 0 11704 400
rect 14952 0 15008 400
rect 18256 0 18312 400
rect 21560 0 21616 400
rect 24864 0 24920 400
rect 28168 0 28224 400
<< obsm2 >>
rect 1638 29570 2938 29600
rect 3054 29570 8930 29600
rect 9046 29570 14922 29600
rect 15038 29570 20914 29600
rect 21030 29570 26906 29600
rect 27022 29570 28714 29600
rect 1638 430 28714 29570
rect 1638 400 1706 430
rect 1822 400 5010 430
rect 5126 400 8314 430
rect 8430 400 11618 430
rect 11734 400 14922 430
rect 15038 400 18226 430
rect 18342 400 21530 430
rect 21646 400 24834 430
rect 24950 400 28138 430
rect 28254 400 28714 430
<< obsm3 >>
rect 2233 1554 28719 28238
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< labels >>
rlabel metal2 s 1736 0 1792 400 6 A[0]
port 1 nsew signal input
rlabel metal2 s 5040 0 5096 400 6 A[1]
port 2 nsew signal input
rlabel metal2 s 8344 0 8400 400 6 A[2]
port 3 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 A[3]
port 4 nsew signal input
rlabel metal2 s 14952 0 15008 400 6 B[0]
port 5 nsew signal input
rlabel metal2 s 18256 0 18312 400 6 B[1]
port 6 nsew signal input
rlabel metal2 s 21560 0 21616 400 6 B[2]
port 7 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 B[3]
port 8 nsew signal input
rlabel metal2 s 2968 29600 3024 30000 6 S[0]
port 9 nsew signal output
rlabel metal2 s 8960 29600 9016 30000 6 S[1]
port 10 nsew signal output
rlabel metal2 s 14952 29600 15008 30000 6 S[2]
port 11 nsew signal output
rlabel metal2 s 20944 29600 21000 30000 6 S[3]
port 12 nsew signal output
rlabel metal2 s 28168 0 28224 400 6 cin
port 13 nsew signal input
rlabel metal2 s 26936 29600 26992 30000 6 cout
port 14 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 15 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 16 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 447842
string GDS_FILE /home/vrushabh/CLA_GF-180/openlane/cla/runs/22_12_05_12_51/results/signoff/cla.magic.gds
string GDS_START 92474
<< end >>

